VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO strongARMLatch
  CLASS CORE ;
  ORIGIN 0.53 -0.27 ;
  FOREIGN strongARMLatch -0.53 0.27 ;
  SIZE 18.07 BY 31.17 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN Voutp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.745 6.69 6.495 6.885 ;
        RECT 6.205 6.665 6.465 6.985 ;
        RECT 4.745 6.665 5.005 6.985 ;
      LAYER li1 ;
        RECT 6.23 7.675 6.4 8.005 ;
        RECT 4.025 17.57 4.22 17.9 ;
        RECT 4.025 17.475 4.195 18.025 ;
        RECT 3.18 5.905 3.365 6.235 ;
        RECT 3.18 5.855 3.35 6.275 ;
        RECT 3.135 9.585 3.315 9.915 ;
        RECT 3.135 9.475 3.305 10.025 ;
      LAYER met1 ;
        RECT 6.205 6.665 6.465 6.985 ;
        RECT 6.2 7.695 6.43 7.985 ;
        RECT 6.225 6.665 6.43 7.985 ;
        RECT 4.745 6.665 5.005 6.985 ;
        RECT 3.995 6.685 5.005 6.96 ;
        RECT 3.975 17.59 4.25 17.88 ;
        RECT 3.935 9.48 4.24 13.735 ;
        RECT 3.995 5.97 4.24 13.735 ;
        RECT 3.975 9.48 4.225 17.88 ;
        RECT 3.51 7.09 4.24 7.465 ;
        RECT 3.165 5.97 4.24 6.15 ;
        RECT 3.115 9.69 4.24 9.855 ;
        RECT 3.165 5.925 3.395 6.215 ;
        RECT 3.115 9.605 3.345 9.895 ;
      LAYER mcon ;
        RECT 3.145 9.665 3.315 9.835 ;
        RECT 3.195 5.985 3.365 6.155 ;
        RECT 4.05 17.65 4.22 17.82 ;
        RECT 6.23 7.755 6.4 7.925 ;
      LAYER via ;
        RECT 4.8 6.75 4.95 6.9 ;
        RECT 6.26 6.75 6.41 6.9 ;
    END
  END Voutp
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 12.245 13.37 12.69 13.92 ;
        RECT 11.325 13.37 11.495 13.92 ;
        RECT 11.295 13.46 11.495 13.79 ;
        RECT 8.13 19.905 8.3 20.455 ;
        RECT 8.125 20.005 8.3 20.335 ;
        RECT 7.365 19.905 7.81 20.455 ;
        RECT 6.945 9.58 7.12 9.91 ;
        RECT 6.945 9.485 7.115 10.035 ;
        RECT 6.18 9.485 6.625 10.035 ;
        RECT 4.515 17.475 4.96 18.025 ;
        RECT 3.595 17.475 3.765 18.025 ;
        RECT 3.555 17.58 3.765 17.91 ;
        RECT 2.675 10.375 3.335 10.645 ;
        RECT 3.055 30.62 3.225 30.95 ;
        RECT 2.705 9.475 2.875 10.025 ;
        RECT 2.695 9.6 2.875 9.93 ;
        RECT 0.425 19.055 0.595 19.605 ;
        RECT 0.42 19.17 0.595 19.5 ;
        RECT -0.34 19.055 0.105 19.605 ;
      LAYER met1 ;
        RECT 10.995 16.505 15.355 17.275 ;
        RECT 14.34 12.795 15.125 17.275 ;
        RECT 12.285 13.23 15.125 13.845 ;
        RECT 12.245 13.37 12.69 13.92 ;
        RECT 7.92 24.695 12.305 25.12 ;
        RECT 10.995 15.125 11.6 25.12 ;
        RECT 10.965 13.21 11.5 15.275 ;
        RECT 7.92 22.38 8.595 30.285 ;
        RECT 8.095 20.025 8.325 20.315 ;
        RECT 8.13 20.025 8.3 20.91 ;
        RECT 8.125 20.595 8.28 30.285 ;
        RECT 7.465 20.775 8.28 21.005 ;
        RECT 2.84 27.24 8.595 28.375 ;
        RECT 7.365 19.905 7.81 20.455 ;
        RECT 7.49 19.905 7.685 21.005 ;
        RECT 5.615 14.96 7.38 15.785 ;
        RECT 6.8 10.25 7.235 15.785 ;
        RECT 6.92 9.6 7.15 9.89 ;
        RECT 6.93 9.6 7.1 15.785 ;
        RECT 2.865 20.945 6.81 21.975 ;
        RECT 5.815 14.96 6.81 21.975 ;
        RECT 6.255 10.795 7.235 11.08 ;
        RECT 6.18 9.485 6.625 10.035 ;
        RECT 6.255 9.485 6.505 11.085 ;
        RECT 4.515 17.585 6.81 17.935 ;
        RECT 4.515 17.475 4.96 18.025 ;
        RECT 2.04 17.6 3.755 17.89 ;
        RECT 2.865 17.385 3.705 30.115 ;
        RECT 2.14 10.375 3.335 10.645 ;
        RECT 3.025 30.64 3.255 30.93 ;
        RECT 3.05 17.385 3.23 30.93 ;
        RECT 2.14 10.365 3.215 10.7 ;
        RECT 2.14 9.62 2.895 9.91 ;
        RECT 2.04 13.86 2.865 20.44 ;
        RECT 2.065 17.385 3.705 20.465 ;
        RECT 0.78 27.33 8.595 28.16 ;
        RECT 2.14 9.605 2.79 20.465 ;
        RECT 0.79 25.63 1.59 28.835 ;
        RECT 0.14 25.535 1.535 25.87 ;
        RECT 0.23 25.63 1.59 26.135 ;
        RECT 0.14 20.69 0.765 25.87 ;
        RECT 0.39 19.19 0.62 19.48 ;
        RECT 0.375 19.255 0.575 26.135 ;
        RECT -0.28 20.075 0.575 20.445 ;
        RECT -0.34 19.055 0.105 19.605 ;
        RECT -0.25 19.055 0.035 20.445 ;
      LAYER mcon ;
        RECT -0.205 19.245 -0.035 19.415 ;
        RECT 0.42 19.25 0.59 19.42 ;
        RECT 2.695 9.68 2.865 9.85 ;
        RECT 2.92 10.425 3.09 10.595 ;
        RECT 3.055 30.7 3.225 30.87 ;
        RECT 3.555 17.66 3.725 17.83 ;
        RECT 4.65 17.665 4.82 17.835 ;
        RECT 6.315 9.675 6.485 9.845 ;
        RECT 6.95 9.66 7.12 9.83 ;
        RECT 7.5 20.095 7.67 20.265 ;
        RECT 8.125 20.085 8.295 20.255 ;
        RECT 11.295 13.54 11.465 13.71 ;
        RECT 12.38 13.56 12.55 13.73 ;
    END
  END VDD
  PIN Voutn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.06 8.52 8.11 8.92 ;
      LAYER li1 ;
        RECT 8.56 20.02 8.735 20.35 ;
        RECT 8.56 19.905 8.73 20.455 ;
        RECT 7.42 6.14 7.59 6.56 ;
        RECT 7.375 9.485 7.545 10.035 ;
        RECT 2.21 7.005 2.38 7.335 ;
      LAYER met1 ;
        RECT 8.46 7.31 9.785 7.58 ;
        RECT 7.345 9.685 8.785 9.845 ;
        RECT 8.515 9.685 8.78 20.26 ;
        RECT 8.535 9.685 8.765 20.33 ;
        RECT 8.465 6.245 8.715 9.845 ;
        RECT 7.39 6.195 8.645 6.43 ;
        RECT 7.915 8.57 8.715 8.88 ;
        RECT 7.845 8.575 8.105 8.895 ;
        RECT 7.39 6.195 7.62 6.5 ;
        RECT 7.345 9.625 7.575 9.915 ;
        RECT 2.18 7.025 2.41 7.315 ;
        RECT 2.135 8.545 2.395 8.865 ;
        RECT 2.115 7.095 2.355 8.84 ;
      LAYER mcon ;
        RECT 2.21 7.085 2.38 7.255 ;
        RECT 7.375 9.685 7.545 9.855 ;
        RECT 7.42 6.27 7.59 6.44 ;
        RECT 8.565 20.1 8.735 20.27 ;
      LAYER via ;
        RECT 2.19 8.63 2.34 8.78 ;
        RECT 7.9 8.66 8.05 8.81 ;
    END
  END Voutn
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 13.08 21.37 17.54 21.955 ;
        RECT 8.515 1.3 17.06 1.88 ;
        RECT 16.265 1.3 16.955 22.06 ;
        RECT 13.51 14.145 16.955 14.855 ;
        RECT 13.465 14.51 16.955 14.83 ;
        RECT 7.17 21.485 17.54 21.765 ;
        RECT 12.005 14.135 12.335 21.765 ;
        RECT 10.315 20.79 10.565 21.765 ;
        RECT 10.265 20.75 10.525 21.07 ;
        RECT 7.17 21.48 9.38 21.77 ;
        RECT 8.95 20.865 9.145 21.77 ;
        RECT 6.355 1.29 9.045 1.65 ;
        RECT 1.6 20.255 7.695 20.485 ;
        RECT 7.17 20.255 7.675 21.84 ;
        RECT 4.505 1.445 6.585 1.82 ;
        RECT 5.225 19 5.43 20.485 ;
        RECT 5.08 18.935 5.34 19.255 ;
        RECT 1.6 20.15 4.995 20.505 ;
        RECT 4.375 1.42 4.635 1.74 ;
        RECT 1.615 19.68 1.82 20.505 ;
        RECT 1.56 19.68 1.82 20 ;
      LAYER li1 ;
        RECT 11.88 14.595 12.05 14.925 ;
        RECT 8.97 20.735 9.14 21.065 ;
        RECT 4 18.92 4.17 19.25 ;
        RECT 3.525 0.98 3.695 1.31 ;
        RECT 1.255 20.23 1.425 20.56 ;
      LAYER met1 ;
        RECT 16.205 23.785 16.85 24.465 ;
        RECT 16.47 21.63 16.73 21.95 ;
        RECT 16.32 21.68 16.695 24.465 ;
        RECT 13.465 14.51 13.725 14.83 ;
        RECT 11.85 14.615 13.655 14.835 ;
        RECT 11.885 14.58 13.725 14.83 ;
        RECT 11.85 14.615 12.08 14.905 ;
        RECT 10.265 20.75 10.525 21.07 ;
        RECT 8.935 20.845 10.525 20.99 ;
        RECT 8.94 20.755 9.17 21.045 ;
        RECT 5.08 18.935 5.34 19.255 ;
        RECT 3.875 19.03 5.34 19.175 ;
        RECT 3.97 18.94 4.2 19.23 ;
        RECT 4.375 1.42 4.635 1.74 ;
        RECT 3.62 1.485 4.635 1.68 ;
        RECT 3.495 1 3.725 1.29 ;
        RECT 3.5 1 3.705 1.64 ;
        RECT 1.06 20.24 1.84 20.49 ;
        RECT 1.56 19.68 1.82 20 ;
        RECT 1.59 19.68 1.79 20.49 ;
        RECT 1.225 20.24 1.455 20.54 ;
      LAYER mcon ;
        RECT 1.255 20.31 1.425 20.48 ;
        RECT 3.525 1.06 3.695 1.23 ;
        RECT 4 19 4.17 19.17 ;
        RECT 8.97 20.815 9.14 20.985 ;
        RECT 11.88 14.675 12.05 14.845 ;
      LAYER via ;
        RECT 1.615 19.765 1.765 19.915 ;
        RECT 4.43 1.505 4.58 1.655 ;
        RECT 5.135 19.02 5.285 19.17 ;
        RECT 10.32 20.835 10.47 20.985 ;
        RECT 13.52 14.595 13.67 14.745 ;
        RECT 16.525 21.715 16.675 21.865 ;
    END
  END clk
  PIN Vinp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.18 4.14 6.35 4.47 ;
      LAYER met1 ;
        RECT 6.15 4.16 6.38 4.45 ;
        RECT 5.545 4.205 6.38 4.445 ;
      LAYER mcon ;
        RECT 6.18 4.22 6.35 4.39 ;
    END
  END Vinp
  PIN Vinn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 3.88 1.635 4.21 ;
      LAYER met1 ;
        RECT 1.435 3.9 1.665 4.19 ;
        RECT 0.445 3.915 1.65 4.225 ;
      LAYER mcon ;
        RECT 1.465 3.96 1.635 4.13 ;
    END
  END Vinn
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 4.835 0.42 5.005 0.84 ;
        RECT 4.825 0.47 5.005 0.8 ;
        RECT 4.15 0.48 4.32 0.81 ;
      LAYER met1 ;
        RECT 4.795 0.49 5.025 0.78 ;
        RECT 4.12 0.53 5.025 0.75 ;
        RECT 4.12 0.5 4.35 0.79 ;
      LAYER mcon ;
        RECT 4.15 0.56 4.32 0.73 ;
        RECT 4.825 0.55 4.995 0.72 ;
    END
  END VSS
  OBS
    LAYER mcon ;
      RECT 11.77 13.555 11.94 13.725 ;
      RECT 7.06 3.355 7.23 3.525 ;
      RECT 6.995 6.275 7.165 6.445 ;
      RECT 6.655 3.31 6.825 3.48 ;
      RECT 5.285 0.54 5.455 0.71 ;
      RECT 2.845 3.23 3.015 3.4 ;
      RECT 2.74 5.99 2.91 6.16 ;
      RECT 2.37 3.22 2.54 3.39 ;
      RECT 0.865 19.255 1.035 19.425 ;
    LAYER met1 ;
      RECT 11.74 13.495 11.97 13.785 ;
      RECT 11.74 4.905 11.915 13.785 ;
      RECT 11.7 4.905 12.015 9.795 ;
      RECT 6.965 6.215 7.195 6.505 ;
      RECT 6.97 5 7.16 6.505 ;
      RECT 6.845 5 8.365 5.23 ;
      RECT 7.78 4.905 12.1 5.17 ;
      RECT 8.135 3.305 8.36 5.23 ;
      RECT 7.03 3.295 7.26 3.585 ;
      RECT 7.03 3.305 8.36 3.505 ;
      RECT 6.625 3.25 6.855 3.54 ;
      RECT 6.655 1.92 6.855 3.54 ;
      RECT 2.365 1.925 2.57 3.475 ;
      RECT 2.34 3.16 2.57 3.45 ;
      RECT 2.38 1.92 6.855 2.125 ;
      RECT 5.295 0.48 5.45 2.125 ;
      RECT 5.255 0.48 5.485 0.77 ;
      RECT 0.835 19.195 1.065 19.485 ;
      RECT 0.86 5.945 1.045 19.485 ;
      RECT 0.85 5.945 1.365 16.96 ;
      RECT 2.71 5.93 2.94 6.22 ;
      RECT 0.85 5.975 2.94 6.145 ;
      RECT 1.92 5.015 2.14 6.145 ;
      RECT 1.92 5.015 3.605 5.24 ;
      RECT 1.92 5.015 3.63 5.23 ;
      RECT 3.46 3.165 3.635 5.115 ;
      RECT 1.93 4.995 3.635 5.115 ;
      RECT 2.755 4.985 3.605 5.24 ;
      RECT 2.815 3.165 3.045 3.46 ;
      RECT 2.815 3.165 3.635 3.395 ;
    LAYER li1 ;
      RECT 11.755 13.37 11.925 13.92 ;
      RECT 11.755 13.475 11.94 13.805 ;
      RECT 7.065 3.2 7.235 3.62 ;
      RECT 7.06 3.275 7.235 3.605 ;
      RECT 6.99 6.14 7.16 6.56 ;
      RECT 6.99 6.195 7.165 6.525 ;
      RECT 6.635 3.2 6.805 3.62 ;
      RECT 6.635 3.23 6.825 3.56 ;
      RECT 5.265 0.42 5.435 0.84 ;
      RECT 5.265 0.46 5.455 0.79 ;
      RECT 2.815 3.095 2.985 3.515 ;
      RECT 2.815 3.15 3.015 3.48 ;
      RECT 2.75 5.855 2.92 6.275 ;
      RECT 2.74 5.91 2.92 6.24 ;
      RECT 2.385 3.095 2.555 3.515 ;
      RECT 2.37 3.14 2.555 3.47 ;
      RECT 0.855 19.055 1.025 19.605 ;
      RECT 0.855 19.175 1.035 19.505 ;
  END
END strongARMLatch

END LIBRARY
